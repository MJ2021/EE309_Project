library ieee;
use ieee.std_logic_1164.all;
use ieee.math_real.all;
use ieee.numeric_std.all;

library work;
use work.components.all;

entity reg_file is
	generic(
		data_length: integer := 16;
		num_reg: integer := 8);
		
	port(
		data_in: in std_logic_vector(data_length-1 downto 0);
		rf_df1, rf_df2, R7_PC: out std_logic_vector(data_length-1 downto 0);
		sel_in, sel_out1, sel_out2: in std_logic_vector(integer(ceil(log2(real(num_reg))))-1 downto 0);
		clk, wr_ena: in std_logic);
		
end entity;

architecture behave of reg_file is
	type data_bus is array(num_reg-1 downto 0) of std_logic_vector(data_length-1 downto 0);
	signal reg_out: data_bus;
	signal ena: std_logic_vector(num_reg-1 downto 0);
	
begin
	
	GEN_REG: 
	for i in 0 to num_reg-1 generate
		REG: reg_process
			generic map(data_length)
			port map(clk => clk, ena => ena(i), 
				Din => data_in, Dout => reg_out(i));
	end generate GEN_REG;
	
	in_decode: process(sel_in, wr_ena)
	begin
		ena <= (others => '0');
		ena(to_integer(unsigned(sel_in))) <= wr_ena;	
	end process;
	
	rf_df1 <= reg_out(to_integer(unsigned(sel_out1)));
	rf_df2 <= reg_out(to_integer(unsigned(sel_out2)));
	R7_PC <= reg_out(num_reg-1);
	
end architecture;